10
10
10
10
10
00
11
11
11
11
11
01
10
10
10
10
00
11
11
11
11
00
